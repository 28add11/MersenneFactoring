`default_nettype none

module square #(
	parameter BITWIDTH=32,
) (
	input wire [BITWIDTH - 1:0] x,
	output reg [BITWIDTH - 1:0] y
);

	
	
endmodule